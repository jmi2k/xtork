typedef struct packed {
	bit[0:3] r;
	bit[0:3] g;
	bit[0:3] b;
} RGB_444;
